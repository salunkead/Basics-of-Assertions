//variable clock delay

/*
##delay 
delay cannot be variable as the delay value must be known before run time.

##[0:lv_data]
in the range operator also variable delay is not possible.

in short,delay values must be constants and it cannot be variables.

what if you want variable delay value?
1. this can be done using local_variable

*/

//Example:-

